// I2C_TOP 
// Author:
// Date: 02/16/2024
// Rev: v0.1
// Description: 
//              v0.1: Inital Version 

module i2c_top();



endmodule